
`timescale 1ns/1ps
module mem_bram #(
    parameter ADDR_WIDTH = 10,		//地址宽度
    parameter DATA_WIDTH = 128		//数据宽度
)(
    input                   clk,   // Clock
    input [ADDR_WIDTH-1:0]  raddr,  // Address
    input [ADDR_WIDTH-1:0]  waddr,  // Address
    input [DATA_WIDTH-1:0]  din,   // Data Input
    input                   we,    // Write Enable
    output [DATA_WIDTH-1:0] dout   // Data Output
); 
    reg [ADDR_WIDTH-1:0] addr_r;  // Address Register
    reg [DATA_WIDTH-1:0] ram [0:(1 << ADDR_WIDTH)-1];
    integer i;
    initial begin
        ram[0][31:0] = 32'd2429146761;
        ram[0][63:32] = 32'd1704984117;
        ram[0][95:64] = 32'd244488320;
        ram[0][127:96] = 32'd2009627834;
        ram[1][31:0] = 32'd1187404859;
        ram[1][63:32] = 32'd1738854148;
        ram[1][95:64] = 32'd120926161;
        ram[1][127:96] = 32'd497144763;
        ram[2][31:0] = 32'd4074274575;
        ram[2][63:32] = 32'd2506404521;
        ram[2][95:64] = 32'd2770097472;
        ram[2][127:96] = 32'd4191856559;
        ram[3][31:0] = 32'd290304978;
        ram[3][63:32] = 32'd3587268486;
        ram[3][95:64] = 32'd2853805329;
        ram[3][127:96] = 32'd618621332;
        ram[4][31:0] = 32'd2339767300;
        ram[4][63:32] = 32'd432400395;
        ram[4][95:64] = 32'd4089621706;
        ram[4][127:96] = 32'd2117409300;
        ram[5][31:0] = 32'd1303944501;
        ram[5][63:32] = 32'd1866610343;
        ram[5][95:64] = 32'd879268720;
        ram[5][127:96] = 32'd291373066;
        ram[6][31:0] = 32'd619906137;
        ram[6][63:32] = 32'd3881438871;
        ram[6][95:64] = 32'd1614175349;
        ram[6][127:96] = 32'd2950000704;
        ram[7][31:0] = 32'd2040897048;
        ram[7][63:32] = 32'd580774497;
        ram[7][95:64] = 32'd4194707533;
        ram[7][127:96] = 32'd1738403846;
        ram[8][31:0] = 32'd695764078;
        ram[8][63:32] = 32'd3369978576;
        ram[8][95:64] = 32'd3084178052;
        ram[8][127:96] = 32'd273674846;
        ram[9][31:0] = 32'd3434138962;
        ram[9][63:32] = 32'd2005231466;
        ram[9][95:64] = 32'd4009161584;
        ram[9][127:96] = 32'd2786481955;
        ram[10][31:0] = 32'd4102836592;
        ram[10][63:32] = 32'd2145959186;
        ram[10][95:64] = 32'd527128804;
        ram[10][127:96] = 32'd3505372607;
        ram[11][31:0] = 32'd3951540326;
        ram[11][63:32] = 32'd1124776585;
        ram[11][95:64] = 32'd1323238552;
        ram[11][127:96] = 32'd2052202513;
        ram[12][31:0] = 32'd4130110526;
        ram[12][63:32] = 32'd1404102730;
        ram[12][95:64] = 32'd2162511413;
        ram[12][127:96] = 32'd2194417863;
        ram[13][31:0] = 32'd1474304506;
        ram[13][63:32] = 32'd1748677916;
        ram[13][95:64] = 32'd2532063245;
        ram[13][127:96] = 32'd2155416609;
        ram[14][31:0] = 32'd2965160517;
        ram[14][63:32] = 32'd2167625309;
        ram[14][95:64] = 32'd3980185017;
        ram[14][127:96] = 32'd587109440;
        ram[15][31:0] = 32'd2464752507;
        ram[15][63:32] = 32'd3065752321;
        ram[15][95:64] = 32'd3712003529;
        ram[15][127:96] = 32'd807961889;
        ram[16][31:0] = 32'd4216388865;
        ram[16][63:32] = 32'd1673314307;
        ram[16][95:64] = 32'd5228628;
        ram[16][127:96] = 32'd283800910;
        ram[17][31:0] = 32'd3879425881;
        ram[17][63:32] = 32'd2408633668;
        ram[17][95:64] = 32'd692439474;
        ram[17][127:96] = 32'd3398690954;
        ram[18][31:0] = 32'd583387573;
        ram[18][63:32] = 32'd1855683855;
        ram[18][95:64] = 32'd1226571034;
        ram[18][127:96] = 32'd1317445743;
        ram[19][31:0] = 32'd2183571412;
        ram[19][63:32] = 32'd1951277074;
        ram[19][95:64] = 32'd3938077862;
        ram[19][127:96] = 32'd3352086201;
        ram[20][31:0] = 32'd3975584697;
        ram[20][63:32] = 32'd1304484359;
        ram[20][95:64] = 32'd2763428529;
        ram[20][127:96] = 32'd1828590022;
        ram[21][31:0] = 32'd1081301073;
        ram[21][63:32] = 32'd725363894;
        ram[21][95:64] = 32'd1595499640;
        ram[21][127:96] = 32'd597900638;
        ram[22][31:0] = 32'd1179514588;
        ram[22][63:32] = 32'd185144842;
        ram[22][95:64] = 32'd43380869;
        ram[22][127:96] = 32'd138001890;
        ram[23][31:0] = 32'd403469968;
        ram[23][63:32] = 32'd563973034;
        ram[23][95:64] = 32'd1435958758;
        ram[23][127:96] = 32'd610452162;
        ram[24][31:0] = 32'd2080744587;
        ram[24][63:32] = 32'd654962339;
        ram[24][95:64] = 32'd3684430035;
        ram[24][127:96] = 32'd1718939551;
        ram[25][31:0] = 32'd3845605637;
        ram[25][63:32] = 32'd669798772;
        ram[25][95:64] = 32'd746597445;
        ram[25][127:96] = 32'd1606109734;
        ram[26][31:0] = 32'd3747696734;
        ram[26][63:32] = 32'd1511183284;
        ram[26][95:64] = 32'd1630641212;
        ram[26][127:96] = 32'd4002934247;
        ram[27][31:0] = 32'd3475654866;
        ram[27][63:32] = 32'd1300879613;
        ram[27][95:64] = 32'd1563193765;
        ram[27][127:96] = 32'd59269632;
        ram[28][31:0] = 32'd26118987;
        ram[28][63:32] = 32'd124869335;
        ram[28][95:64] = 32'd2347304629;
        ram[28][127:96] = 32'd2227853741;
        ram[29][31:0] = 32'd3242481180;
        ram[29][63:32] = 32'd3928372404;
        ram[29][95:64] = 32'd2838500611;
        ram[29][127:96] = 32'd2525938397;
        ram[30][31:0] = 32'd3491273784;
        ram[30][63:32] = 32'd539709361;
        ram[30][95:64] = 32'd3741684855;
        ram[30][127:96] = 32'd2458661410;
        ram[31][31:0] = 32'd3922973245;
        ram[31][63:32] = 32'd1835274807;
        ram[31][95:64] = 32'd4195730453;
        ram[31][127:96] = 32'd598873427;
        ram[32][31:0] = 32'd3391204038;
        ram[32][63:32] = 32'd652071928;
        ram[32][95:64] = 32'd246684452;
        ram[32][127:96] = 32'd1010540666;
        ram[33][31:0] = 32'd3352808087;
        ram[33][63:32] = 32'd2182795532;
        ram[33][95:64] = 32'd2143987429;
        ram[33][127:96] = 32'd2176215843;
        ram[34][31:0] = 32'd3446836288;
        ram[34][63:32] = 32'd2464351703;
        ram[34][95:64] = 32'd1330454173;
        ram[34][127:96] = 32'd3027351263;
        ram[35][31:0] = 32'd3314446855;
        ram[35][63:32] = 32'd1108123326;
        ram[35][95:64] = 32'd3762198714;
        ram[35][127:96] = 32'd1862437858;
        ram[36][31:0] = 32'd1832364570;
        ram[36][63:32] = 32'd2945026917;
        ram[36][95:64] = 32'd3958907471;
        ram[36][127:96] = 32'd3396137010;
        ram[37][31:0] = 32'd3092460397;
        ram[37][63:32] = 32'd3842519337;
        ram[37][95:64] = 32'd2726814038;
        ram[37][127:96] = 32'd1136502393;
        ram[38][31:0] = 32'd800774714;
        ram[38][63:32] = 32'd3239039963;
        ram[38][95:64] = 32'd3022540257;
        ram[38][127:96] = 32'd3939648809;
        ram[39][31:0] = 32'd2004451240;
        ram[39][63:32] = 32'd98365346;
        ram[39][95:64] = 32'd2430407245;
        ram[39][127:96] = 32'd3077284633;
        ram[40][31:0] = 32'd2802001540;
        ram[40][63:32] = 32'd260760954;
        ram[40][95:64] = 32'd760186910;
        ram[40][127:96] = 32'd2417096706;
        ram[41][31:0] = 32'd3847429411;
        ram[41][63:32] = 32'd309152437;
        ram[41][95:64] = 32'd1567391663;
        ram[41][127:96] = 32'd4201079425;
        ram[42][31:0] = 32'd244697080;
        ram[42][63:32] = 32'd49778203;
        ram[42][95:64] = 32'd900511560;
        ram[42][127:96] = 32'd1827178944;
        ram[43][31:0] = 32'd2706684257;
        ram[43][63:32] = 32'd1739717906;
        ram[43][95:64] = 32'd3406369137;
        ram[43][127:96] = 32'd1951074742;
        ram[44][31:0] = 32'd3605693122;
        ram[44][63:32] = 32'd934387763;
        ram[44][95:64] = 32'd1390194371;
        ram[44][127:96] = 32'd4169806564;
        ram[45][31:0] = 32'd2888358889;
        ram[45][63:32] = 32'd485480945;
        ram[45][95:64] = 32'd407882722;
        ram[45][127:96] = 32'd1700753432;
        ram[46][31:0] = 32'd4125218622;
        ram[46][63:32] = 32'd3591529659;
        ram[46][95:64] = 32'd621023615;
        ram[46][127:96] = 32'd329709741;
        ram[47][31:0] = 32'd3828919794;
        ram[47][63:32] = 32'd2152553771;
        ram[47][95:64] = 32'd2871768144;
        ram[47][127:96] = 32'd211975995;
        ram[48][31:0] = 32'd3438095621;
        ram[48][63:32] = 32'd1908158991;
        ram[48][95:64] = 32'd3455513250;
        ram[48][127:96] = 32'd3242935053;
        ram[49][31:0] = 32'd3889204301;
        ram[49][63:32] = 32'd3675913621;
        ram[49][95:64] = 32'd400801465;
        ram[49][127:96] = 32'd3233870748;
        ram[50][31:0] = 32'd3223549335;
        ram[50][63:32] = 32'd2012336102;
        ram[50][95:64] = 32'd631181234;
        ram[50][127:96] = 32'd827013616;
        ram[51][31:0] = 32'd218891852;
        ram[51][63:32] = 32'd540360476;
        ram[51][95:64] = 32'd2946247101;
        ram[51][127:96] = 32'd689273551;
        ram[52][31:0] = 32'd1843892378;
        ram[52][63:32] = 32'd76413089;
        ram[52][95:64] = 32'd788019105;
        ram[52][127:96] = 32'd3948687695;
        ram[53][31:0] = 32'd3169469609;
        ram[53][63:32] = 32'd2763846381;
        ram[53][95:64] = 32'd3563881117;
        ram[53][127:96] = 32'd2441226058;
        ram[54][31:0] = 32'd313568208;
        ram[54][63:32] = 32'd2658004276;
        ram[54][95:64] = 32'd3295815568;
        ram[54][127:96] = 32'd1970268263;
        ram[55][31:0] = 32'd3319839920;
        ram[55][63:32] = 32'd2679756236;
        ram[55][95:64] = 32'd2498690093;
        ram[55][127:96] = 32'd3261764772;
        ram[56][31:0] = 32'd4068853398;
        ram[56][63:32] = 32'd1364845516;
        ram[56][95:64] = 32'd3088560151;
        ram[56][127:96] = 32'd4109066461;
        ram[57][31:0] = 32'd2455014083;
        ram[57][63:32] = 32'd2383148880;
        ram[57][95:64] = 32'd2673908551;
        ram[57][127:96] = 32'd3679121765;
        ram[58][31:0] = 32'd3657253458;
        ram[58][63:32] = 32'd894914896;
        ram[58][95:64] = 32'd2569948806;
        ram[58][127:96] = 32'd2173127971;
        ram[59][31:0] = 32'd1629491404;
        ram[59][63:32] = 32'd2163671273;
        ram[59][95:64] = 32'd1309914105;
        ram[59][127:96] = 32'd2680540905;
        ram[60][31:0] = 32'd4111033551;
        ram[60][63:32] = 32'd738113948;
        ram[60][95:64] = 32'd2340774178;
        ram[60][127:96] = 32'd309132402;
        ram[61][31:0] = 32'd3986444448;
        ram[61][63:32] = 32'd3305055470;
        ram[61][95:64] = 32'd2440705799;
        ram[61][127:96] = 32'd873071231;
        ram[62][31:0] = 32'd1851737756;
        ram[62][63:32] = 32'd4121500431;
        ram[62][95:64] = 32'd1892908102;
        ram[62][127:96] = 32'd402216612;
        ram[63][31:0] = 32'd2678663684;
        ram[63][63:32] = 32'd1046892784;
        ram[63][95:64] = 32'd893686890;
        ram[63][127:96] = 32'd738701221;
        ram[64][31:0] = 32'd104124540;
        ram[64][63:32] = 32'd2272834637;
        ram[64][95:64] = 32'd2183547082;
        ram[64][127:96] = 32'd3199409289;
        ram[65][31:0] = 32'd3784376997;
        ram[65][63:32] = 32'd3435254937;
        ram[65][95:64] = 32'd2953460781;
        ram[65][127:96] = 32'd1168259603;
        ram[66][31:0] = 32'd3017312274;
        ram[66][63:32] = 32'd4232753553;
        ram[66][95:64] = 32'd4193755358;
        ram[66][127:96] = 32'd2420869187;
        ram[67][31:0] = 32'd2644833872;
        ram[67][63:32] = 32'd2018394395;
        ram[67][95:64] = 32'd245427783;
        ram[67][127:96] = 32'd4226387963;
        ram[68][31:0] = 32'd1785668236;
        ram[68][63:32] = 32'd3957578884;
        ram[68][95:64] = 32'd3297475855;
        ram[68][127:96] = 32'd3441919684;
        ram[69][31:0] = 32'd151084863;
        ram[69][63:32] = 32'd1313409944;
        ram[69][95:64] = 32'd3951155712;
        ram[69][127:96] = 32'd2152272633;
        ram[70][31:0] = 32'd1318904363;
        ram[70][63:32] = 32'd2803364487;
        ram[70][95:64] = 32'd3250739478;
        ram[70][127:96] = 32'd1573656911;
        ram[71][31:0] = 32'd2237941646;
        ram[71][63:32] = 32'd1224676552;
        ram[71][95:64] = 32'd1413268032;
        ram[71][127:96] = 32'd1630502931;
        ram[72][31:0] = 32'd2933858888;
        ram[72][63:32] = 32'd2358155133;
        ram[72][95:64] = 32'd1764399317;
        ram[72][127:96] = 32'd2014839919;
        ram[73][31:0] = 32'd149615558;
        ram[73][63:32] = 32'd880389596;
        ram[73][95:64] = 32'd2673885267;
        ram[73][127:96] = 32'd1453477040;
        ram[74][31:0] = 32'd72603561;
        ram[74][63:32] = 32'd1556985237;
        ram[74][95:64] = 32'd189733476;
        ram[74][127:96] = 32'd1004966428;
        ram[75][31:0] = 32'd1786211448;
        ram[75][63:32] = 32'd2613515428;
        ram[75][95:64] = 32'd3250392161;
        ram[75][127:96] = 32'd4095352313;
        ram[76][31:0] = 32'd3750445638;
        ram[76][63:32] = 32'd129216807;
        ram[76][95:64] = 32'd480752041;
        ram[76][127:96] = 32'd4030103948;
        ram[77][31:0] = 32'd2797128928;
        ram[77][63:32] = 32'd1328657515;
        ram[77][95:64] = 32'd3828155493;
        ram[77][127:96] = 32'd3422864683;
        ram[78][31:0] = 32'd2136184510;
        ram[78][63:32] = 32'd3975800125;
        ram[78][95:64] = 32'd1771827745;
        ram[78][127:96] = 32'd1180062760;
        ram[79][31:0] = 32'd1714277137;
        ram[79][63:32] = 32'd613544344;
        ram[79][95:64] = 32'd1356147939;
        ram[79][127:96] = 32'd180363106;
        ram[80][31:0] = 32'd4010594226;
        ram[80][63:32] = 32'd2130141956;
        ram[80][95:64] = 32'd2434467256;
        ram[80][127:96] = 32'd1823069783;
        ram[81][31:0] = 32'd4124680673;
        ram[81][63:32] = 32'd1292476535;
        ram[81][95:64] = 32'd3245783896;
        ram[81][127:96] = 32'd4021375997;
        ram[82][31:0] = 32'd4211559137;
        ram[82][63:32] = 32'd508970632;
        ram[82][95:64] = 32'd2871069657;
        ram[82][127:96] = 32'd1391651160;
        ram[83][31:0] = 32'd1631465858;
        ram[83][63:32] = 32'd3777587601;
        ram[83][95:64] = 32'd2560750633;
        ram[83][127:96] = 32'd3132902255;
        ram[84][31:0] = 32'd535597245;
        ram[84][63:32] = 32'd2803068549;
        ram[84][95:64] = 32'd1957293410;
        ram[84][127:96] = 32'd1615140309;
        ram[85][31:0] = 32'd3854321255;
        ram[85][63:32] = 32'd3105826626;
        ram[85][95:64] = 32'd148146141;
        ram[85][127:96] = 32'd3938949624;
        ram[86][31:0] = 32'd477263003;
        ram[86][63:32] = 32'd1569155127;
        ram[86][95:64] = 32'd4150117994;
        ram[86][127:96] = 32'd4057955162;
        ram[87][31:0] = 32'd3314453200;
        ram[87][63:32] = 32'd992540281;
        ram[87][95:64] = 32'd1842231339;
        ram[87][127:96] = 32'd435348931;
        ram[88][31:0] = 32'd2176341776;
        ram[88][63:32] = 32'd2052389658;
        ram[88][95:64] = 32'd369923590;
        ram[88][127:96] = 32'd2603783369;
        ram[89][31:0] = 32'd3608961784;
        ram[89][63:32] = 32'd1704996566;
        ram[89][95:64] = 32'd3479819972;
        ram[89][127:96] = 32'd309287193;
        ram[90][31:0] = 32'd1414751202;
        ram[90][63:32] = 32'd2280030852;
        ram[90][95:64] = 32'd883421312;
        ram[90][127:96] = 32'd3362159751;
        ram[91][31:0] = 32'd4091092656;
        ram[91][63:32] = 32'd1876322875;
        ram[91][95:64] = 32'd2904869292;
        ram[91][127:96] = 32'd1478079112;
        ram[92][31:0] = 32'd1594529834;
        ram[92][63:32] = 32'd1912926533;
        ram[92][95:64] = 32'd3118834818;
        ram[92][127:96] = 32'd1688419579;
        ram[93][31:0] = 32'd3823632809;
        ram[93][63:32] = 32'd3237219661;
        ram[93][95:64] = 32'd149363693;
        ram[93][127:96] = 32'd2093158352;
        ram[94][31:0] = 32'd736569085;
        ram[94][63:32] = 32'd1111968953;
        ram[94][95:64] = 32'd4089108044;
        ram[94][127:96] = 32'd2445988135;
        ram[95][31:0] = 32'd2614266083;
        ram[95][63:32] = 32'd3380814185;
        ram[95][95:64] = 32'd2573507917;
        ram[95][127:96] = 32'd2516549088;
        ram[96][31:0] = 32'd739005625;
        ram[96][63:32] = 32'd698224158;
        ram[96][95:64] = 32'd1877039969;
        ram[96][127:96] = 32'd140765230;
        ram[97][31:0] = 32'd640328259;
        ram[97][63:32] = 32'd2090137532;
        ram[97][95:64] = 32'd2928158067;
        ram[97][127:96] = 32'd1779555079;
        ram[98][31:0] = 32'd10599762;
        ram[98][63:32] = 32'd1215078312;
        ram[98][95:64] = 32'd2899126994;
        ram[98][127:96] = 32'd4037953191;
        ram[99][31:0] = 32'd150757965;
        ram[99][63:32] = 32'd3740595799;
        ram[99][95:64] = 32'd1885338136;
        ram[99][127:96] = 32'd798523023;
        ram[100][31:0] = 32'd12061985;
        ram[100][63:32] = 32'd1367308988;
        ram[100][95:64] = 32'd3328109157;
        ram[100][127:96] = 32'd1931821484;
        ram[101][31:0] = 32'd1720976526;
        ram[101][63:32] = 32'd3263563325;
        ram[101][95:64] = 32'd380969902;
        ram[101][127:96] = 32'd3124378955;
        ram[102][31:0] = 32'd3784952382;
        ram[102][63:32] = 32'd829691805;
        ram[102][95:64] = 32'd1292454337;
        ram[102][127:96] = 32'd1053791089;
        ram[103][31:0] = 32'd1038301027;
        ram[103][63:32] = 32'd2856665508;
        ram[103][95:64] = 32'd1136158832;
        ram[103][127:96] = 32'd268942874;
        ram[104][31:0] = 32'd2315947450;
        ram[104][63:32] = 32'd2168180925;
        ram[104][95:64] = 32'd1834403807;
        ram[104][127:96] = 32'd3511401386;
        ram[105][31:0] = 32'd2422752708;
        ram[105][63:32] = 32'd257964552;
        ram[105][95:64] = 32'd962672775;
        ram[105][127:96] = 32'd3728980285;
        ram[106][31:0] = 32'd974442485;
        ram[106][63:32] = 32'd3494559305;
        ram[106][95:64] = 32'd3544872180;
        ram[106][127:96] = 32'd2561035456;
        ram[107][31:0] = 32'd3571198896;
        ram[107][63:32] = 32'd3277805322;
        ram[107][95:64] = 32'd1822620302;
        ram[107][127:96] = 32'd1854590995;
        ram[108][31:0] = 32'd3691339593;
        ram[108][63:32] = 32'd2768242345;
        ram[108][95:64] = 32'd3036540911;
        ram[108][127:96] = 32'd1857893028;
        ram[109][31:0] = 32'd1804759271;
        ram[109][63:32] = 32'd446220078;
        ram[109][95:64] = 32'd943277004;
        ram[109][127:96] = 32'd1055579969;
        ram[110][31:0] = 32'd867078260;
        ram[110][63:32] = 32'd700898576;
        ram[110][95:64] = 32'd2814803870;
        ram[110][127:96] = 32'd1114978954;
        ram[111][31:0] = 32'd2972090766;
        ram[111][63:32] = 32'd1931819170;
        ram[111][95:64] = 32'd421789546;
        ram[111][127:96] = 32'd1470049012;
        ram[112][31:0] = 32'd3836817188;
        ram[112][63:32] = 32'd1938256718;
        ram[112][95:64] = 32'd2419356892;
        ram[112][127:96] = 32'd869464472;
        ram[113][31:0] = 32'd1443069133;
        ram[113][63:32] = 32'd3913516686;
        ram[113][95:64] = 32'd3918291114;
        ram[113][127:96] = 32'd131669732;
        ram[114][31:0] = 32'd2655493248;
        ram[114][63:32] = 32'd2493953492;
        ram[114][95:64] = 32'd2786993620;
        ram[114][127:96] = 32'd576195236;
        ram[115][31:0] = 32'd1397313540;
        ram[115][63:32] = 32'd3896793757;
        ram[115][95:64] = 32'd954874650;
        ram[115][127:96] = 32'd2623477901;
        ram[116][31:0] = 32'd2727706364;
        ram[116][63:32] = 32'd2741905062;
        ram[116][95:64] = 32'd3459645207;
        ram[116][127:96] = 32'd4019651710;
        ram[117][31:0] = 32'd3992930714;
        ram[117][63:32] = 32'd1664670904;
        ram[117][95:64] = 32'd43804014;
        ram[117][127:96] = 32'd3733821095;
        ram[118][31:0] = 32'd463884868;
        ram[118][63:32] = 32'd1293966191;
        ram[118][95:64] = 32'd95842768;
        ram[118][127:96] = 32'd2268014519;
        ram[119][31:0] = 32'd3560019982;
        ram[119][63:32] = 32'd3221152013;
        ram[119][95:64] = 32'd3294322927;
        ram[119][127:96] = 32'd2603322669;
        ram[120][31:0] = 32'd338748893;
        ram[120][63:32] = 32'd3104519648;
        ram[120][95:64] = 32'd2959940318;
        ram[120][127:96] = 32'd2078207425;
        ram[121][31:0] = 32'd1372237211;
        ram[121][63:32] = 32'd3869014208;
        ram[121][95:64] = 32'd1136344694;
        ram[121][127:96] = 32'd397506953;
        ram[122][31:0] = 32'd3725295247;
        ram[122][63:32] = 32'd2421545610;
        ram[122][95:64] = 32'd3475954419;
        ram[122][127:96] = 32'd3079598917;
        ram[123][31:0] = 32'd712901222;
        ram[123][63:32] = 32'd712725379;
        ram[123][95:64] = 32'd602403619;
        ram[123][127:96] = 32'd3266638749;
        ram[124][31:0] = 32'd822810503;
        ram[124][63:32] = 32'd1711199328;
        ram[124][95:64] = 32'd3738045385;
        ram[124][127:96] = 32'd3460457963;
        ram[125][31:0] = 32'd2119686540;
        ram[125][63:32] = 32'd2870347926;
        ram[125][95:64] = 32'd2391045745;
        ram[125][127:96] = 32'd2345310091;
        ram[126][31:0] = 32'd2260143172;
        ram[126][63:32] = 32'd413069247;
        ram[126][95:64] = 32'd998035363;
        ram[126][127:96] = 32'd724258612;
        ram[127][31:0] = 32'd3350070891;
        ram[127][63:32] = 32'd2006610656;
        ram[127][95:64] = 32'd4129103904;
        ram[127][127:96] = 32'd1421325492;
        ram[128][31:0] = 32'd3788029954;
        ram[128][63:32] = 32'd1638524148;
        ram[128][95:64] = 32'd1160262532;
        ram[128][127:96] = 32'd2354318472;
        ram[129][31:0] = 32'd173393108;
        ram[129][63:32] = 32'd2393872258;
        ram[129][95:64] = 32'd1538424755;
        ram[129][127:96] = 32'd705002716;
        ram[130][31:0] = 32'd3688177324;
        ram[130][63:32] = 32'd1306264201;
        ram[130][95:64] = 32'd2366573361;
        ram[130][127:96] = 32'd1659053730;
        ram[131][31:0] = 32'd2535488802;
        ram[131][63:32] = 32'd1473714708;
        ram[131][95:64] = 32'd3009779400;
        ram[131][127:96] = 32'd3043177996;
        ram[132][31:0] = 32'd1208414750;
        ram[132][63:32] = 32'd1896802361;
        ram[132][95:64] = 32'd1192716121;
        ram[132][127:96] = 32'd1530930906;
        ram[133][31:0] = 32'd1329842884;
        ram[133][63:32] = 32'd3593280808;
        ram[133][95:64] = 32'd1623632665;
        ram[133][127:96] = 32'd1728180162;
        ram[134][31:0] = 32'd2953848538;
        ram[134][63:32] = 32'd367782055;
        ram[134][95:64] = 32'd2395926350;
        ram[134][127:96] = 32'd3897175329;
        ram[135][31:0] = 32'd2220496832;
        ram[135][63:32] = 32'd1920105602;
        ram[135][95:64] = 32'd3693452330;
        ram[135][127:96] = 32'd1985053232;
        ram[136][31:0] = 32'd118999468;
        ram[136][63:32] = 32'd1749290836;
        ram[136][95:64] = 32'd717909476;
        ram[136][127:96] = 32'd1656097789;
        ram[137][31:0] = 32'd3975122350;
        ram[137][63:32] = 32'd2127589844;
        ram[137][95:64] = 32'd2320911093;
        ram[137][127:96] = 32'd604963152;
        ram[138][31:0] = 32'd1286678884;
        ram[138][63:32] = 32'd1687299562;
        ram[138][95:64] = 32'd3923557028;
        ram[138][127:96] = 32'd2248499919;
        ram[139][31:0] = 32'd2939472687;
        ram[139][63:32] = 32'd985122537;
        ram[139][95:64] = 32'd3808977718;
        ram[139][127:96] = 32'd839457297;
        ram[140][31:0] = 32'd2158590197;
        ram[140][63:32] = 32'd2792998988;
        ram[140][95:64] = 32'd1942238216;
        ram[140][127:96] = 32'd3656355596;
        ram[141][31:0] = 32'd1073823995;
        ram[141][63:32] = 32'd1483039500;
        ram[141][95:64] = 32'd3645197110;
        ram[141][127:96] = 32'd3156642332;
        ram[142][31:0] = 32'd148205842;
        ram[142][63:32] = 32'd4106722886;
        ram[142][95:64] = 32'd1424901878;
        ram[142][127:96] = 32'd4031278286;
        ram[143][31:0] = 32'd894425430;
        ram[143][63:32] = 32'd1409403198;
        ram[143][95:64] = 32'd2569024098;
        ram[143][127:96] = 32'd1100236442;
        ram[144][31:0] = 32'd2445404047;
        ram[144][63:32] = 32'd513421463;
        ram[144][95:64] = 32'd2894820147;
        ram[144][127:96] = 32'd3224225652;
        ram[145][31:0] = 32'd1239202064;
        ram[145][63:32] = 32'd2716519087;
        ram[145][95:64] = 32'd1383356002;
        ram[145][127:96] = 32'd2544097139;
        ram[146][31:0] = 32'd2050130973;
        ram[146][63:32] = 32'd791050687;
        ram[146][95:64] = 32'd3389351130;
        ram[146][127:96] = 32'd3912203569;
        ram[147][31:0] = 32'd2997617910;
        ram[147][63:32] = 32'd788551438;
        ram[147][95:64] = 32'd763136854;
        ram[147][127:96] = 32'd2476460923;
        ram[148][31:0] = 32'd3656952568;
        ram[148][63:32] = 32'd767211102;
        ram[148][95:64] = 32'd2232370504;
        ram[148][127:96] = 32'd2295987580;
        ram[149][31:0] = 32'd3890943431;
        ram[149][63:32] = 32'd4054056191;
        ram[149][95:64] = 32'd133191090;
        ram[149][127:96] = 32'd1504995887;
        ram[150][31:0] = 32'd1736910815;
        ram[150][63:32] = 32'd1528966083;
        ram[150][95:64] = 32'd2985258556;
        ram[150][127:96] = 32'd1521945037;
        ram[151][31:0] = 32'd2635934467;
        ram[151][63:32] = 32'd3385414901;
        ram[151][95:64] = 32'd3060791752;
        ram[151][127:96] = 32'd3129915412;
        ram[152][31:0] = 32'd4173859586;
        ram[152][63:32] = 32'd2651952637;
        ram[152][95:64] = 32'd2655954426;
        ram[152][127:96] = 32'd507597236;
        ram[153][31:0] = 32'd3082247360;
        ram[153][63:32] = 32'd98227944;
        ram[153][95:64] = 32'd2818354787;
        ram[153][127:96] = 32'd3553517321;
        ram[154][31:0] = 32'd1763094828;
        ram[154][63:32] = 32'd15484412;
        ram[154][95:64] = 32'd2989005313;
        ram[154][127:96] = 32'd2093912685;
        ram[155][31:0] = 32'd23215832;
        ram[155][63:32] = 32'd2767751789;
        ram[155][95:64] = 32'd3415325110;
        ram[155][127:96] = 32'd2296683503;
        ram[156][31:0] = 32'd50566768;
        ram[156][63:32] = 32'd1546441285;
        ram[156][95:64] = 32'd1317854929;
        ram[156][127:96] = 32'd2223197704;
        ram[157][31:0] = 32'd228558971;
        ram[157][63:32] = 32'd1662750713;
        ram[157][95:64] = 32'd732867767;
        ram[157][127:96] = 32'd2020367395;
        ram[158][31:0] = 32'd2717021060;
        ram[158][63:32] = 32'd3017373220;
        ram[158][95:64] = 32'd2429702712;
        ram[158][127:96] = 32'd1607332002;
        ram[159][31:0] = 32'd3849721588;
        ram[159][63:32] = 32'd3517993239;
        ram[159][95:64] = 32'd4136659456;
        ram[159][127:96] = 32'd86901798;
        ram[160][31:0] = 32'd3316842311;
        ram[160][63:32] = 32'd741175375;
        ram[160][95:64] = 32'd3003817392;
        ram[160][127:96] = 32'd1955210064;
        ram[161][31:0] = 32'd2998446653;
        ram[161][63:32] = 32'd1474811439;
        ram[161][95:64] = 32'd1560612810;
        ram[161][127:96] = 32'd360683726;
        ram[162][31:0] = 32'd2360713956;
        ram[162][63:32] = 32'd3974071841;
        ram[162][95:64] = 32'd4203221935;
        ram[162][127:96] = 32'd3706032235;
        ram[163][31:0] = 32'd3888780918;
        ram[163][63:32] = 32'd923572889;
        ram[163][95:64] = 32'd3014930614;
        ram[163][127:96] = 32'd2201370237;
        ram[164][31:0] = 32'd2492457321;
        ram[164][63:32] = 32'd576451002;
        ram[164][95:64] = 32'd2306672925;
        ram[164][127:96] = 32'd4136402978;
        ram[165][31:0] = 32'd2587946543;
        ram[165][63:32] = 32'd1404351648;
        ram[165][95:64] = 32'd4126887004;
        ram[165][127:96] = 32'd3355262986;
        ram[166][31:0] = 32'd1318050398;
        ram[166][63:32] = 32'd1327055600;
        ram[166][95:64] = 32'd3537140051;
        ram[166][127:96] = 32'd1268036190;
        ram[167][31:0] = 32'd1499949566;
        ram[167][63:32] = 32'd3091727096;
        ram[167][95:64] = 32'd2901628700;
        ram[167][127:96] = 32'd3009182528;
        ram[168][31:0] = 32'd442134545;
        ram[168][63:32] = 32'd3204904385;
        ram[168][95:64] = 32'd824316215;
        ram[168][127:96] = 32'd2709261325;
        ram[169][31:0] = 32'd1104785019;
        ram[169][63:32] = 32'd1594126675;
        ram[169][95:64] = 32'd4257693411;
        ram[169][127:96] = 32'd3806169552;
        ram[170][31:0] = 32'd111880350;
        ram[170][63:32] = 32'd1236016341;
        ram[170][95:64] = 32'd3033798570;
        ram[170][127:96] = 32'd3097106317;
        ram[171][31:0] = 32'd1377128895;
        ram[171][63:32] = 32'd992539895;
        ram[171][95:64] = 32'd626729407;
        ram[171][127:96] = 32'd2332656559;
        ram[172][31:0] = 32'd903539134;
        ram[172][63:32] = 32'd2479435461;
        ram[172][95:64] = 32'd1799699601;
        ram[172][127:96] = 32'd1926809194;
        ram[173][31:0] = 32'd3393115954;
        ram[173][63:32] = 32'd1755618517;
        ram[173][95:64] = 32'd1783902209;
        ram[173][127:96] = 32'd4120276502;
        ram[174][31:0] = 32'd1053390424;
        ram[174][63:32] = 32'd150212881;
        ram[174][95:64] = 32'd259042086;
        ram[174][127:96] = 32'd3824988992;
        ram[175][31:0] = 32'd2431932061;
        ram[175][63:32] = 32'd835744670;
        ram[175][95:64] = 32'd3588029089;
        ram[175][127:96] = 32'd1255659046;
        ram[176][31:0] = 32'd998116682;
        ram[176][63:32] = 32'd503495629;
        ram[176][95:64] = 32'd1013806716;
        ram[176][127:96] = 32'd1113132010;
        ram[177][31:0] = 32'd3884518045;
        ram[177][63:32] = 32'd3130440955;
        ram[177][95:64] = 32'd3654683160;
        ram[177][127:96] = 32'd1104666845;
        ram[178][31:0] = 32'd3993640537;
        ram[178][63:32] = 32'd3877347980;
        ram[178][95:64] = 32'd1793666688;
        ram[178][127:96] = 32'd701885885;
        ram[179][31:0] = 32'd2594539979;
        ram[179][63:32] = 32'd4165932764;
        ram[179][95:64] = 32'd2871267844;
        ram[179][127:96] = 32'd3591465327;
        ram[180][31:0] = 32'd2657030068;
        ram[180][63:32] = 32'd662721243;
        ram[180][95:64] = 32'd4264062206;
        ram[180][127:96] = 32'd2035228107;
        ram[181][31:0] = 32'd3488346519;
        ram[181][63:32] = 32'd4023969800;
        ram[181][95:64] = 32'd1456997450;
        ram[181][127:96] = 32'd2168181148;
        ram[182][31:0] = 32'd716320088;
        ram[182][63:32] = 32'd3068713767;
        ram[182][95:64] = 32'd3458672318;
        ram[182][127:96] = 32'd1618801135;
        ram[183][31:0] = 32'd1195362064;
        ram[183][63:32] = 32'd844566830;
        ram[183][95:64] = 32'd1357887344;
        ram[183][127:96] = 32'd4218761319;
        ram[184][31:0] = 32'd914072280;
        ram[184][63:32] = 32'd565879052;
        ram[184][95:64] = 32'd3739241179;
        ram[184][127:96] = 32'd2457990130;
        ram[185][31:0] = 32'd2567066062;
        ram[185][63:32] = 32'd2013379092;
        ram[185][95:64] = 32'd546339758;
        ram[185][127:96] = 32'd2720583043;
        ram[186][31:0] = 32'd4202166401;
        ram[186][63:32] = 32'd3734504505;
        ram[186][95:64] = 32'd2402779610;
        ram[186][127:96] = 32'd4029219969;
        ram[187][31:0] = 32'd1620627030;
        ram[187][63:32] = 32'd428043726;
        ram[187][95:64] = 32'd632044382;
        ram[187][127:96] = 32'd500787216;
        ram[188][31:0] = 32'd3981528151;
        ram[188][63:32] = 32'd3199516579;
        ram[188][95:64] = 32'd733598019;
        ram[188][127:96] = 32'd3037275798;
        ram[189][31:0] = 32'd943611231;
        ram[189][63:32] = 32'd2785722476;
        ram[189][95:64] = 32'd848987015;
        ram[189][127:96] = 32'd290937831;
        ram[190][31:0] = 32'd2415159896;
        ram[190][63:32] = 32'd1930378489;
        ram[190][95:64] = 32'd2315924990;
        ram[190][127:96] = 32'd3670633852;
        ram[191][31:0] = 32'd3480601920;
        ram[191][63:32] = 32'd549136353;
        ram[191][95:64] = 32'd1936387940;
        ram[191][127:96] = 32'd1779844196;
        ram[192][31:0] = 32'd3269737958;
        ram[192][63:32] = 32'd855063859;
        ram[192][95:64] = 32'd2728342669;
        ram[192][127:96] = 32'd2140434203;
        ram[193][31:0] = 32'd2174708313;
        ram[193][63:32] = 32'd3204087429;
        ram[193][95:64] = 32'd773021249;
        ram[193][127:96] = 32'd193689677;
        ram[194][31:0] = 32'd2103915868;
        ram[194][63:32] = 32'd3351668101;
        ram[194][95:64] = 32'd1485151742;
        ram[194][127:96] = 32'd25730636;
        ram[195][31:0] = 32'd3449249766;
        ram[195][63:32] = 32'd2618963896;
        ram[195][95:64] = 32'd1895287559;
        ram[195][127:96] = 32'd840459236;
        ram[196][31:0] = 32'd2409029183;
        ram[196][63:32] = 32'd1730244568;
        ram[196][95:64] = 32'd4210699665;
        ram[196][127:96] = 32'd3191758865;
        ram[197][31:0] = 32'd3817033739;
        ram[197][63:32] = 32'd484067223;
        ram[197][95:64] = 32'd1938234177;
        ram[197][127:96] = 32'd3456993164;
        ram[198][31:0] = 32'd3388575783;
        ram[198][63:32] = 32'd1843129498;
        ram[198][95:64] = 32'd350349391;
        ram[198][127:96] = 32'd1540072738;
        ram[199][31:0] = 32'd1292528924;
        ram[199][63:32] = 32'd3703456760;
        ram[199][95:64] = 32'd2831706730;
        ram[199][127:96] = 32'd1361996462;
        ram[200][31:0] = 32'd2684303926;
        ram[200][63:32] = 32'd2873799072;
        ram[200][95:64] = 32'd3491622919;
        ram[200][127:96] = 32'd3660731959;
        ram[201][31:0] = 32'd2619582498;
        ram[201][63:32] = 32'd341095953;
        ram[201][95:64] = 32'd3109763568;
        ram[201][127:96] = 32'd619472320;
        ram[202][31:0] = 32'd3811340329;
        ram[202][63:32] = 32'd3174497928;
        ram[202][95:64] = 32'd848075204;
        ram[202][127:96] = 32'd1022680166;
        ram[203][31:0] = 32'd732597252;
        ram[203][63:32] = 32'd2469749640;
        ram[203][95:64] = 32'd3911919694;
        ram[203][127:96] = 32'd4204391240;
        ram[204][31:0] = 32'd3714792815;
        ram[204][63:32] = 32'd3647515413;
        ram[204][95:64] = 32'd3263948359;
        ram[204][127:96] = 32'd2910897927;
        ram[205][31:0] = 32'd2587666766;
        ram[205][63:32] = 32'd3918583867;
        ram[205][95:64] = 32'd3241601505;
        ram[205][127:96] = 32'd3228310104;
        ram[206][31:0] = 32'd1705558585;
        ram[206][63:32] = 32'd3901277367;
        ram[206][95:64] = 32'd1621627116;
        ram[206][127:96] = 32'd4087048189;
        ram[207][31:0] = 32'd3346872234;
        ram[207][63:32] = 32'd275433189;
        ram[207][95:64] = 32'd3958563769;
        ram[207][127:96] = 32'd3088253311;
        ram[208][31:0] = 32'd2891161115;
        ram[208][63:32] = 32'd1793456890;
        ram[208][95:64] = 32'd3031697508;
        ram[208][127:96] = 32'd1220150061;
        ram[209][31:0] = 32'd319479514;
        ram[209][63:32] = 32'd2699943669;
        ram[209][95:64] = 32'd2155428742;
        ram[209][127:96] = 32'd2174987116;
        ram[210][31:0] = 32'd403783328;
        ram[210][63:32] = 32'd846659615;
        ram[210][95:64] = 32'd3536331538;
        ram[210][127:96] = 32'd1817785861;
        ram[211][31:0] = 32'd1900608026;
        ram[211][63:32] = 32'd2737759682;
        ram[211][95:64] = 32'd3605947957;
        ram[211][127:96] = 32'd2773855860;
        ram[212][31:0] = 32'd2760016426;
        ram[212][63:32] = 32'd644666857;
        ram[212][95:64] = 32'd3810045984;
        ram[212][127:96] = 32'd1633202550;
        ram[213][31:0] = 32'd3434666825;
        ram[213][63:32] = 32'd564835311;
        ram[213][95:64] = 32'd2378975131;
        ram[213][127:96] = 32'd3981959618;
        ram[214][31:0] = 32'd821321256;
        ram[214][63:32] = 32'd54187291;
        ram[214][95:64] = 32'd1198553052;
        ram[214][127:96] = 32'd3073653273;
        ram[215][31:0] = 32'd3552320581;
        ram[215][63:32] = 32'd469402357;
        ram[215][95:64] = 32'd3411959600;
        ram[215][127:96] = 32'd3900994997;
        ram[216][31:0] = 32'd2448373667;
        ram[216][63:32] = 32'd3891425040;
        ram[216][95:64] = 32'd366355984;
        ram[216][127:96] = 32'd566958024;
        ram[217][31:0] = 32'd1380517056;
        ram[217][63:32] = 32'd2551007028;
        ram[217][95:64] = 32'd612456591;
        ram[217][127:96] = 32'd1653013973;
        ram[218][31:0] = 32'd44098560;
        ram[218][63:32] = 32'd2989369719;
        ram[218][95:64] = 32'd3038300328;
        ram[218][127:96] = 32'd931550812;
        ram[219][31:0] = 32'd2137203319;
        ram[219][63:32] = 32'd1774453158;
        ram[219][95:64] = 32'd1205002421;
        ram[219][127:96] = 32'd2912634867;
        ram[220][31:0] = 32'd2614693622;
        ram[220][63:32] = 32'd1107971482;
        ram[220][95:64] = 32'd809342124;
        ram[220][127:96] = 32'd997878904;
        ram[221][31:0] = 32'd665306548;
        ram[221][63:32] = 32'd1599653647;
        ram[221][95:64] = 32'd2973579849;
        ram[221][127:96] = 32'd2450826475;
        ram[222][31:0] = 32'd3501273103;
        ram[222][63:32] = 32'd858761786;
        ram[222][95:64] = 32'd3932332099;
        ram[222][127:96] = 32'd1541522239;
        ram[223][31:0] = 32'd1705100511;
        ram[223][63:32] = 32'd2641599984;
        ram[223][95:64] = 32'd1045852187;
        ram[223][127:96] = 32'd119509833;
        ram[224][31:0] = 32'd298321624;
        ram[224][63:32] = 32'd2281912767;
        ram[224][95:64] = 32'd262579741;
        ram[224][127:96] = 32'd3207744075;
        ram[225][31:0] = 32'd3651982289;
        ram[225][63:32] = 32'd1575034248;
        ram[225][95:64] = 32'd910704321;
        ram[225][127:96] = 32'd242028171;
        ram[226][31:0] = 32'd2673042208;
        ram[226][63:32] = 32'd3640324962;
        ram[226][95:64] = 32'd774256557;
        ram[226][127:96] = 32'd901261549;
        ram[227][31:0] = 32'd2319053902;
        ram[227][63:32] = 32'd1140222346;
        ram[227][95:64] = 32'd885454967;
        ram[227][127:96] = 32'd1201879819;
        ram[228][31:0] = 32'd624833006;
        ram[228][63:32] = 32'd3108154670;
        ram[228][95:64] = 32'd4156785633;
        ram[228][127:96] = 32'd1563133648;
        ram[229][31:0] = 32'd755342212;
        ram[229][63:32] = 32'd4071938350;
        ram[229][95:64] = 32'd3107554339;
        ram[229][127:96] = 32'd2511923435;
        ram[230][31:0] = 32'd3915123610;
        ram[230][63:32] = 32'd3532290497;
        ram[230][95:64] = 32'd181860439;
        ram[230][127:96] = 32'd1705989553;
        ram[231][31:0] = 32'd2793887872;
        ram[231][63:32] = 32'd1313195782;
        ram[231][95:64] = 32'd2215204705;
        ram[231][127:96] = 32'd877988174;
        ram[232][31:0] = 32'd3715639018;
        ram[232][63:32] = 32'd1467497009;
        ram[232][95:64] = 32'd1729249679;
        ram[232][127:96] = 32'd1776715744;
        ram[233][31:0] = 32'd360085129;
        ram[233][63:32] = 32'd893437629;
        ram[233][95:64] = 32'd392045396;
        ram[233][127:96] = 32'd2632191667;
        ram[234][31:0] = 32'd3408512394;
        ram[234][63:32] = 32'd3663858100;
        ram[234][95:64] = 32'd3969264942;
        ram[234][127:96] = 32'd4240778167;
        ram[235][31:0] = 32'd338549878;
        ram[235][63:32] = 32'd2633217852;
        ram[235][95:64] = 32'd2811349348;
        ram[235][127:96] = 32'd3145560359;
        ram[236][31:0] = 32'd1901157862;
        ram[236][63:32] = 32'd2616613166;
        ram[236][95:64] = 32'd4251511846;
        ram[236][127:96] = 32'd2403214353;
        ram[237][31:0] = 32'd990983367;
        ram[237][63:32] = 32'd525044368;
        ram[237][95:64] = 32'd2680314078;
        ram[237][127:96] = 32'd2339532244;
        ram[238][31:0] = 32'd4040559479;
        ram[238][63:32] = 32'd2421064545;
        ram[238][95:64] = 32'd920008339;
        ram[238][127:96] = 32'd3697128996;
        ram[239][31:0] = 32'd922515263;
        ram[239][63:32] = 32'd2955972127;
        ram[239][95:64] = 32'd1131678623;
        ram[239][127:96] = 32'd3011059689;
        ram[240][31:0] = 32'd813414639;
        ram[240][63:32] = 32'd2648618923;
        ram[240][95:64] = 32'd3660914740;
        ram[240][127:96] = 32'd3778906056;
        ram[241][31:0] = 32'd1676243570;
        ram[241][63:32] = 32'd533232901;
        ram[241][95:64] = 32'd168242151;
        ram[241][127:96] = 32'd2540554632;
        ram[242][31:0] = 32'd759450314;
        ram[242][63:32] = 32'd4246657183;
        ram[242][95:64] = 32'd1523162636;
        ram[242][127:96] = 32'd1160760996;
        ram[243][31:0] = 32'd764522856;
        ram[243][63:32] = 32'd1572552106;
        ram[243][95:64] = 32'd3026688618;
        ram[243][127:96] = 32'd902628290;
        ram[244][31:0] = 32'd882564056;
        ram[244][63:32] = 32'd275231142;
        ram[244][95:64] = 32'd452232048;
        ram[244][127:96] = 32'd2852800281;
        ram[245][31:0] = 32'd2034359482;
        ram[245][63:32] = 32'd3011134919;
        ram[245][95:64] = 32'd4040828699;
        ram[245][127:96] = 32'd1211923792;
        ram[246][31:0] = 32'd1238370014;
        ram[246][63:32] = 32'd1224700992;
        ram[246][95:64] = 32'd1388652941;
        ram[246][127:96] = 32'd3353173506;
        ram[247][31:0] = 32'd2478676154;
        ram[247][63:32] = 32'd3635546882;
        ram[247][95:64] = 32'd718330319;
        ram[247][127:96] = 32'd461026114;
        ram[248][31:0] = 32'd2125549255;
        ram[248][63:32] = 32'd1857244546;
        ram[248][95:64] = 32'd2089204886;
        ram[248][127:96] = 32'd3226654615;
        ram[249][31:0] = 32'd3922015050;
        ram[249][63:32] = 32'd1759334156;
        ram[249][95:64] = 32'd143133281;
        ram[249][127:96] = 32'd3093736890;
        ram[250][31:0] = 32'd2546864569;
        ram[250][63:32] = 32'd326676280;
        ram[250][95:64] = 32'd3643312403;
        ram[250][127:96] = 32'd1542999208;
        ram[251][31:0] = 32'd2413861351;
        ram[251][63:32] = 32'd3126585085;
        ram[251][95:64] = 32'd2573864613;
        ram[251][127:96] = 32'd166563627;
        ram[252][31:0] = 32'd4215858546;
        ram[252][63:32] = 32'd1316389492;
        ram[252][95:64] = 32'd3511528593;
        ram[252][127:96] = 32'd70628960;
        ram[253][31:0] = 32'd1486798971;
        ram[253][63:32] = 32'd1056707852;
        ram[253][95:64] = 32'd414447015;
        ram[253][127:96] = 32'd4068782698;
        ram[254][31:0] = 32'd379732789;
        ram[254][63:32] = 32'd3652225397;
        ram[254][95:64] = 32'd2984861369;
        ram[254][127:96] = 32'd4093193534;
        ram[255][31:0] = 32'd1171431187;
        ram[255][63:32] = 32'd3036274148;
        ram[255][95:64] = 32'd657762763;
        ram[255][127:96] = 32'd2095860060;

    end
    always @(posedge clk) begin
        addr_r <= raddr;
        if(we) ram[waddr] <= din;
    end
    assign dout = ram[addr_r]; 

endmodule
